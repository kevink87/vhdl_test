library ieee;

use ieee.std_logic_1164.all;

entity wrapper is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity wrapper;

architecture RTL of wrapper is
	
begin

end architecture RTL;
